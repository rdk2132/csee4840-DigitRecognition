module MAC (input clk, reset
            input signed [15:0] A, B
            output signed [15:0] output)
//Control circuitry for CNN
module CNN_ctrl();

endmodule